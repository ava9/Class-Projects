library verilog;
use verilog.vl_types.all;
entity Decoder is
    generic(
        RTYPE           : vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi1, Hi1);
        OTHER           : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        BRANCH          : vl_logic_vector(1 downto 0) := (Hi1, Hi0);
        ADD             : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        SUB             : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        \SRA\           : vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi0);
        \SRL\           : vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        \SLL\           : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        \AND\           : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi1);
        \OR\            : vl_logic_vector(2 downto 0) := (Hi1, Hi1, Hi0);
        LB              : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi0);
        PSB             : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi0, Hi0);
        ADDI            : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi0, Hi1);
        ANDI            : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi1, Hi0);
        ORI             : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi1, Hi1);
        BEQ             : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        BNE             : vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        BGEZ            : vl_logic_vector(1 downto 0) := (Hi1, Hi0);
        BLTZ            : vl_logic_vector(1 downto 0) := (Hi1, Hi1)
    );
    port(
        INSTR           : in     vl_logic_vector(15 downto 0);
        DR              : out    vl_logic_vector(2 downto 0);
        SA              : out    vl_logic_vector(2 downto 0);
        SB              : out    vl_logic_vector(2 downto 0);
        IMMO            : out    vl_logic_vector(5 downto 0);
        MB              : out    vl_logic;
        FS              : out    vl_logic_vector(2 downto 0);
        MD              : out    vl_logic;
        LD              : out    vl_logic;
        MW              : out    vl_logic;
        HALT            : out    vl_logic;
        BS              : out    vl_logic_vector(2 downto 0);
        OFF             : out    vl_logic_vector(5 downto 0)
    );
    attribute RTYPE_mti_vect_attrib : integer;
    attribute RTYPE_mti_vect_attrib of RTYPE : constant is 15;
    attribute OTHER_mti_vect_attrib : integer;
    attribute OTHER_mti_vect_attrib of OTHER : constant is 0;
    attribute BRANCH_mti_vect_attrib : integer;
    attribute BRANCH_mti_vect_attrib of BRANCH : constant is 2;
    attribute ADD_mti_vect_attrib : integer;
    attribute ADD_mti_vect_attrib of ADD : constant is 0;
    attribute SUB_mti_vect_attrib : integer;
    attribute SUB_mti_vect_attrib of SUB : constant is 1;
    attribute \SRA\\_mti_vect_attrib\ : integer;
    attribute \SRA\\_mti_vect_attrib\ of \SRA\ : constant is 2;
    attribute \SRL\\_mti_vect_attrib\ : integer;
    attribute \SRL\\_mti_vect_attrib\ of \SRL\ : constant is 3;
    attribute \SLL\\_mti_vect_attrib\ : integer;
    attribute \SLL\\_mti_vect_attrib\ of \SLL\ : constant is 4;
    attribute \AND\\_mti_vect_attrib\ : integer;
    attribute \AND\\_mti_vect_attrib\ of \AND\ : constant is 5;
    attribute \OR\\_mti_vect_attrib\ : integer;
    attribute \OR\\_mti_vect_attrib\ of \OR\ : constant is 6;
    attribute LB_mti_vect_attrib : integer;
    attribute LB_mti_vect_attrib of LB : constant is 2;
    attribute PSB_mti_vect_attrib : integer;
    attribute PSB_mti_vect_attrib of PSB : constant is 4;
    attribute ADDI_mti_vect_attrib : integer;
    attribute ADDI_mti_vect_attrib of ADDI : constant is 5;
    attribute ANDI_mti_vect_attrib : integer;
    attribute ANDI_mti_vect_attrib of ANDI : constant is 6;
    attribute ORI_mti_vect_attrib : integer;
    attribute ORI_mti_vect_attrib of ORI : constant is 7;
    attribute BEQ_mti_vect_attrib : integer;
    attribute BEQ_mti_vect_attrib of BEQ : constant is 0;
    attribute BNE_mti_vect_attrib : integer;
    attribute BNE_mti_vect_attrib of BNE : constant is 1;
    attribute BGEZ_mti_vect_attrib : integer;
    attribute BGEZ_mti_vect_attrib of BGEZ : constant is 2;
    attribute BLTZ_mti_vect_attrib : integer;
    attribute BLTZ_mti_vect_attrib of BLTZ : constant is 3;
end Decoder;
