module lab5iram2A(CLK, RESET, ADDR, Q);
  input         CLK;
  input         RESET;
  input  [7:0]  ADDR;
  output [15:0] Q;

  reg    [15:0] mem[0:127]; // instruction memory with 16 bit entries

  wire   [6:0]  saddr;
  integer       i;


  assign saddr = ADDR[7:1];
  assign Q = mem[saddr];

  always @(posedge CLK) begin
    if(RESET) begin
      mem[0]   <= 16'b1111010010010001;   // SUB  R2, R2, R2
      mem[1]   <= 16'b1111001001001001;   // SUB  R1, R1, R1
      mem[2]   <= 16'b0101010010111111;   // ADDI R2, R2, -1
      mem[3]   <= 16'b0100010001000000;   // SB   R1, 0(R2)
      mem[4]   <= 16'b0101001001000001;   // ADDI R1, R1, 1
      mem[5]   <= 16'b0100010001000000;   // SB   R1, 0(R2)
      mem[6]   <= 16'b0101001001000001;   // ADDI R1, R1, 1
      mem[7]   <= 16'b0100010001000000;   // SB   R1, 0(R2)
      mem[8]   <= 16'b0000000000000001;   // HALT
      mem[9]   <= 16'b0101001001000001;   // ADDI R1, R1, 1
      mem[10]  <= 16'b0100010001000000;   // SB   R1, 0(R2)
      mem[11]  <= 16'b0000000000000001;   // HALT
      mem[12]  <= 16'b0101001001000001;   // ADDI R1, R1, 1
      mem[13]  <= 16'b0100010001000000;   // SB   R1, 0(R2)
      mem[14]  <= 16'b0101001001000001;   // ADDI R1, R1, 1
      mem[15]  <= 16'b0100010001000000;   // SB   R1, 0(R2)
      mem[16]  <= 16'b0000000000000001;   // HALT
      mem[17]  <= 16'b1111011011011001;   // SUB  R3, R3, R3
      mem[18]  <= 16'b0101011011000001;   // ADDI R3, R3, 1
      mem[19]  <= 16'b1111001011001000;   // ADD  R1, R1, R3
      mem[20]  <= 16'b0100010001000000;   // SB   R1, 0(R2)
      mem[21]  <= 16'b1111011001001110;   // OR   R1, R3, R1
      mem[22]  <= 16'b0100010001000000;   // SB   R1, 0(R2)
      mem[23]  <= 16'b0000000000000001;   // HALT
      mem[24]  <= 16'b0101011001000000;   // ADDI R1, R3, 0
      mem[25]  <= 16'b1111001000001100;   // SLL  R1, R1
      mem[26]  <= 16'b1111001000001100;   // SLL  R1, R1
      mem[27]  <= 16'b1111001000001100;   // SLL  R1, R1
      mem[28]  <= 16'b0100010001000000;   // SB   R1, 0(R2)
      mem[29]  <= 16'b0111001001000001;   // ORI  R1, R1, 1
      mem[30]  <= 16'b0100010001000000;   // SB   R1, 0(R2)
      mem[31]  <= 16'b0100011001000000;   // SB   R1, 0(R3)
      mem[32]  <= 16'b1111011011011001;   // SUB  R3, R3, R3
      mem[33]  <= 16'b0010011011000001;   // LB   R3, 1(R3)
      mem[34]  <= 16'b0101011001000001;   // ADDI R1, R3, 1
      mem[35]  <= 16'b0100010001000000;   // SB   R1, 0(R2)
      mem[36]  <= 16'b1111001000001100;   // SLL  R1, R1
      mem[37]  <= 16'b1111001000001100;   // SLL  R1, R1
      mem[38]  <= 16'b0101001001101110;   // ADDI R1, R1, -18
      mem[39]  <= 16'b1111001000001011;   // SRL  R1, R1
      mem[40]  <= 16'b0100010001000000;   // SB   R1, 0(R2)
      mem[41]  <= 16'b0000000000000001;   // HALT
      mem[42]  <= 16'b0000000000000000;   // NOP
      mem[43]  <= 16'b0000000000000000;   // NOP
      mem[44]  <= 16'b0101001001000001;   // ADDI R1, R1, 1
      mem[45]  <= 16'b1111010000010010;   // SRA  R2, R2
      mem[46]  <= 16'b0100010001000000;   // SB   R1, 0(R2)
      mem[47]  <= 16'b0110010100011010;   // ANDI R4, R2, 26
      mem[48]  <= 16'b1111100000100010;   // SRA  R4, R4
      mem[49]  <= 16'b0100010100000000;   // SB   R4, 0(R2)
      mem[50]  <= 16'b0000000000000001;   // HALT
      mem[51]  <= 16'b0101011111111110;   // ADDI R7, R3, -2
      mem[52]  <= 16'b1111111010000101;   // AND  R0, R7, R2
      mem[53]  <= 16'b1111000000101000;   // ADD  R5, R0, R0
      mem[54]  <= 16'b0100010101000000;   // SB   R5, 0(R2)

      for(i = 55; i < 128; i = i + 1) begin
        mem[i] <= 16'b0000000000000000;
      end
    end
  end

endmodule
